library verilog;
use verilog.vl_types.all;
entity phaseDecoder_vlg_vec_tst is
end phaseDecoder_vlg_vec_tst;
