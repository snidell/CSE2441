library verilog;
use verilog.vl_types.all;
entity \Lab4DE1-2\ is
    port(
        Sum             : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        Cin             : in     vl_logic;
        Carryout        : out    vl_logic
    );
end \Lab4DE1-2\;
