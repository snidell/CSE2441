library verilog;
use verilog.vl_types.all;
entity opDecoder_vlg_vec_tst is
end opDecoder_vlg_vec_tst;
