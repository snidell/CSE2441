library verilog;
use verilog.vl_types.all;
entity accController_vlg_vec_tst is
end accController_vlg_vec_tst;
