library verilog;
use verilog.vl_types.all;
entity Lab4DE2_vlg_vec_tst is
end Lab4DE2_vlg_vec_tst;
