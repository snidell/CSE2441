library verilog;
use verilog.vl_types.all;
entity homeworkProb_vlg_vec_tst is
end homeworkProb_vlg_vec_tst;
