library verilog;
use verilog.vl_types.all;
entity Lab3AdderSubtractor_vlg_vec_tst is
end Lab3AdderSubtractor_vlg_vec_tst;
