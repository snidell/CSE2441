library verilog;
use verilog.vl_types.all;
entity Lab2Adder_vlg_vec_tst is
end Lab2Adder_vlg_vec_tst;
