library verilog;
use verilog.vl_types.all;
entity slide10pointone_vlg_vec_tst is
end slide10pointone_vlg_vec_tst;
