library verilog;
use verilog.vl_types.all;
entity FourBitTwistedRingCounter_vlg_vec_tst is
end FourBitTwistedRingCounter_vlg_vec_tst;
