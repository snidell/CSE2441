library verilog;
use verilog.vl_types.all;
entity Lab4DE2_vlg_check_tst is
    port(
        Carryout        : in     vl_logic;
        Sum             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab4DE2_vlg_check_tst;
