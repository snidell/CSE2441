library verilog;
use verilog.vl_types.all;
entity RippleAdder_vlg_vec_tst is
end RippleAdder_vlg_vec_tst;
