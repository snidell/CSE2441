library verilog;
use verilog.vl_types.all;
entity slide10pointone_vlg_check_tst is
    port(
        Z1              : in     vl_logic;
        Z2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end slide10pointone_vlg_check_tst;
