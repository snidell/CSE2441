library verilog;
use verilog.vl_types.all;
entity Lab2Adder_vlg_check_tst is
    port(
        P               : in     vl_logic;
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab2Adder_vlg_check_tst;
